`timescale 1ns/1ps
//`define USE_MEM

module memory
  #(
    parameter MEM_FILE = "/home/suyash/git/urisc/example/a.out"
    )(
      input 			   clk,
      
      input [gc::WORD_SIZE - 1:0] 	   add1,
      input [gc::WORD_SIZE - 1:0] 	   dataIn1,
      input 			   write1,
      output reg [gc::WORD_SIZE - 1:0] dataOut1,
      
      input [gc::WORD_SIZE - 1:0] 	   add2,
      input [gc::WORD_SIZE - 1:0] 	   dataIn2,
      input 			   write2,
      output reg [gc::WORD_SIZE - 1:0] dataOut2
      );
   
   (* ram_style = "block" *) reg [gc::WORD_SIZE-1:0] mem [gc::MEM_SIZE - 1:0];

   integer 			   fileID;
   reg [gc::WORD_SIZE-1:0] word;
   integer r, f;

`ifndef USE_MEM
   initial begin
       mem[0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[1] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
       mem[2] = 64'b0000000000000000000000000000000000000000000000000000000000000010;
       mem[3] = 64'b0000000000000000000000000000000000000000000000000000000000000011;
       mem[4] = 64'b0000000000000000000000000000000000000000000000000000000000000100;
       mem[5] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[6] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[7] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[8] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[9] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[10] = 64'b0000000000000000000010110000000000000000001100000000000000000011;
       mem[11] = 64'b0000000000000000000011000000000000000000001100000000000010000001;
       mem[12] = 64'b0000000000000000000011010000000000000000010000000000000000000100;
       mem[13] = 64'b0000000000000000000011100000000000000000010000000000000000000011;
       mem[14] = 64'b0000000000000000000010100000000000000000000000000000000000000000;
       mem[15] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[16] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[17] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[18] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[19] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[20] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[21] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[22] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[23] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[24] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[25] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[26] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[27] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[28] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[29] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[30] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[31] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[32] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[33] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[34] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[35] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[36] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[37] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[38] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[39] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[40] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[41] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[42] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[43] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[44] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[45] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[46] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[47] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[48] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[49] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[50] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[51] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[52] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[53] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[54] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[55] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[56] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[57] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[58] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[59] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[60] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[61] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[62] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[63] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[64] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[65] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[66] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[67] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[68] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[69] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[70] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[71] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[72] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[73] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[74] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[75] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[76] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[77] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[78] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[79] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[80] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[81] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[82] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[83] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[84] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[85] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[86] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[87] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[88] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[89] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[90] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[91] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[92] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[93] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[94] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[95] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[96] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[97] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[98] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[99] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[100] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[101] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[102] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[103] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[104] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[105] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[106] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[107] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[108] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
       mem[109] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
   end
`endif

   always @(posedge clk) begin
   #1
       if (write1) begin
	   mem[add1] <= dataIn1;
       end else begin
	   dataOut1 <= mem[add1];
       end
   end
   
   always @(posedge clk) begin
   #1
       if (write2) begin
	   mem[add2] <= dataIn2;
       end else begin
	   dataOut2 <= mem[add2];
       end
   end
endmodule // memory
