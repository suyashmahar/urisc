`ifndef __VGA_CONSTANTS_VERILOG_HEADER__
`define __VGA_CONSTANTS_VERILOG_HEADER__

parameter SCREEN_HEIGHT = 480;
parameter SCREEN_WIDTH = 640;

parameter LINE_WIDTH = 80, LINE_COUNT = 30;
parameter CHAR_WIDTH = 8, CHAR_HEIGHT = 16;

parameter ROM_SIZE = 128*CHAR_HEIGHT;
parameter ASCII_SIZE = 8;

parameter CHARS_VERT = SCREEN_HEIGHT/CHAR_HEIGHT;
parameter CHARS_HORZ = SCREEN_WIDTH/CHAR_WIDTH;
`endif //  `ifndef __VGA_CONSTANTS_VERILOG_HEADER__
