/*
 * Contains globals package for project wide variables 
 */

package gc; // Global Constants
   parameter WORD_SIZE = 16;
   parameter MEM_SIZE = 1024;
endpackage : gc// globals
   
