`ifndef __URISC_URISC_SV_HEADER__
 `define __URISC_URISC_SV_HEADER__

 `include "cFunctions.svh"
import gc::*;
import utils::*;

`endif      
